`include "i2c_base_test.sv"
`include "i2c_simple_test.sv" 
`include "i2c_address_test.sv"
`include "i2c_spec_addr_reg_order_no_adc_test.sv"
`include "i2c_spec_addr_reg_order_adc_test.sv"
`include "i2c_invalid_address_test.sv"
`include "i2c_invalid_regs_test.sv"
`include "i2c_invalid_adc_write_test.sv"
`include "i2c_all_in_one_test.sv"
`include "i2c_adc_test.sv"
`include "i2c_testing_test.sv"
